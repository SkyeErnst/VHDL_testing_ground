library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity RegAdderTest_TB is
end entity RegAdderTest_TB;